//=====================================================================
// Project: 4 core MESI cache design
// File Name: test_lib.svh
// Description: Base test class and list of tests
// Designers: Venky & Suru
//=====================================================================
//TODO: add your testcase files in here
`include "base_test.sv"
`include "read_miss_icache.sv"
//`include "randomised.sv"
`include "cache_data_miss_read.sv"
`include "cache_data_hit_read.sv"
`include "cache_data_miss_write.sv"
`include "cache_data_hit_write.sv"
`include "cache_inst_hit_read.sv"
